0
0 0 0 0 0 h 2 T 3 B 5 H
0 0 0 0 0 h 2 T
0 0 0 0 0 h 1 B 5 H
0 0 0 0 0 h 6 B 7 B
