0
20 24 20 19 19 r 38 43 47 55 h 25 T 30 B 37 T
20 20 20 20 20 r 48 56 64 h 32 H 44 B
20 20 20 22 20 r 24 33 41 50 h 16 H 40 B
20 20 20 20 20 r 27 32 h 20 H 27 H
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9 
